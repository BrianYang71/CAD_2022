module top(in1, in2, in3, out1);
  input [3:0] in1, in2, in3;
  output [3:0] out1;
  wire [3:0] in1, in2, in3;
  wire [3:0] out1;
  wire csa_tree_ADD_TC_OP_groupi_n_0, csa_tree_ADD_TC_OP_groupi_n_1, csa_tree_ADD_TC_OP_groupi_n_2, csa_tree_ADD_TC_OP_groupi_n_3, csa_tree_ADD_TC_OP_groupi_n_4, csa_tree_ADD_TC_OP_groupi_n_5, csa_tree_ADD_TC_OP_groupi_n_6, csa_tree_ADD_TC_OP_groupi_n_7;
  wire csa_tree_ADD_TC_OP_groupi_n_8, csa_tree_ADD_TC_OP_groupi_n_9, csa_tree_ADD_TC_OP_groupi_n_10, csa_tree_ADD_TC_OP_groupi_n_11, csa_tree_ADD_TC_OP_groupi_n_12, csa_tree_ADD_TC_OP_groupi_n_13, csa_tree_ADD_TC_OP_groupi_n_14, csa_tree_ADD_TC_OP_groupi_n_15;
  wire csa_tree_ADD_TC_OP_groupi_n_16, csa_tree_ADD_TC_OP_groupi_n_17, csa_tree_ADD_TC_OP_groupi_n_18, csa_tree_ADD_TC_OP_groupi_n_19, csa_tree_ADD_TC_OP_groupi_n_20, csa_tree_ADD_TC_OP_groupi_n_21, csa_tree_ADD_TC_OP_groupi_n_22, csa_tree_ADD_TC_OP_groupi_n_23;
  wire csa_tree_ADD_TC_OP_groupi_n_24, csa_tree_ADD_TC_OP_groupi_n_25, csa_tree_ADD_TC_OP_groupi_n_26, csa_tree_ADD_TC_OP_groupi_n_27, csa_tree_ADD_TC_OP_groupi_n_28, csa_tree_ADD_TC_OP_groupi_n_29, csa_tree_ADD_TC_OP_groupi_n_30, csa_tree_ADD_TC_OP_groupi_n_31;
  wire csa_tree_ADD_TC_OP_groupi_n_32, csa_tree_ADD_TC_OP_groupi_n_33, csa_tree_ADD_TC_OP_groupi_n_34, csa_tree_ADD_TC_OP_groupi_n_35, csa_tree_ADD_TC_OP_groupi_n_36, csa_tree_ADD_TC_OP_groupi_n_37, csa_tree_ADD_TC_OP_groupi_n_39, csa_tree_ADD_TC_OP_groupi_n_40;
  wire csa_tree_ADD_TC_OP_groupi_n_41, csa_tree_ADD_TC_OP_groupi_n_42, csa_tree_ADD_TC_OP_groupi_n_43, csa_tree_ADD_TC_OP_groupi_n_44, csa_tree_ADD_TC_OP_groupi_n_45, csa_tree_ADD_TC_OP_groupi_n_46, csa_tree_ADD_TC_OP_groupi_n_47, csa_tree_ADD_TC_OP_groupi_n_48;
  wire csa_tree_ADD_TC_OP_groupi_n_49, csa_tree_ADD_TC_OP_groupi_n_50, csa_tree_ADD_TC_OP_groupi_n_51, csa_tree_ADD_TC_OP_groupi_n_53, csa_tree_ADD_TC_OP_groupi_n_54, csa_tree_ADD_TC_OP_groupi_n_55;
  assign out1[3] = ~(csa_tree_ADD_TC_OP_groupi_n_54  ^ csa_tree_ADD_TC_OP_groupi_n_55 );
  assign out1[2] = ~(csa_tree_ADD_TC_OP_groupi_n_48  ^ csa_tree_ADD_TC_OP_groupi_n_0 );
  assign csa_tree_ADD_TC_OP_groupi_n_55 = ~(csa_tree_ADD_TC_OP_groupi_n_46  ^ csa_tree_ADD_TC_OP_groupi_n_51 );
  assign csa_tree_ADD_TC_OP_groupi_n_54 = ~(csa_tree_ADD_TC_OP_groupi_n_50  | csa_tree_ADD_TC_OP_groupi_n_53 );
  assign csa_tree_ADD_TC_OP_groupi_n_53 = ~(csa_tree_ADD_TC_OP_groupi_n_48  | csa_tree_ADD_TC_OP_groupi_n_49 );
  assign out1[1] = ~(csa_tree_ADD_TC_OP_groupi_n_31  ^ csa_tree_ADD_TC_OP_groupi_n_45 );
  assign csa_tree_ADD_TC_OP_groupi_n_51 = ~(csa_tree_ADD_TC_OP_groupi_n_42  ^ csa_tree_ADD_TC_OP_groupi_n_43 );
  assign csa_tree_ADD_TC_OP_groupi_n_50 = csa_tree_ADD_TC_OP_groupi_n_30  & csa_tree_ADD_TC_OP_groupi_n_44 ;
  assign csa_tree_ADD_TC_OP_groupi_n_49 = ~(csa_tree_ADD_TC_OP_groupi_n_30  | csa_tree_ADD_TC_OP_groupi_n_44 );
  assign csa_tree_ADD_TC_OP_groupi_n_48 = csa_tree_ADD_TC_OP_groupi_n_39  & csa_tree_ADD_TC_OP_groupi_n_47 ;
  assign csa_tree_ADD_TC_OP_groupi_n_47 = csa_tree_ADD_TC_OP_groupi_n_31  | csa_tree_ADD_TC_OP_groupi_n_41 ;
  assign csa_tree_ADD_TC_OP_groupi_n_46 = ~(csa_tree_ADD_TC_OP_groupi_n_28  | csa_tree_ADD_TC_OP_groupi_n_40 );
  assign csa_tree_ADD_TC_OP_groupi_n_45 = ~(csa_tree_ADD_TC_OP_groupi_n_21  ^ csa_tree_ADD_TC_OP_groupi_n_36 );
  assign csa_tree_ADD_TC_OP_groupi_n_44 = ~(csa_tree_ADD_TC_OP_groupi_n_37  ^ csa_tree_ADD_TC_OP_groupi_n_33 );
  assign csa_tree_ADD_TC_OP_groupi_n_43 = ~(csa_tree_ADD_TC_OP_groupi_n_22  ^ csa_tree_ADD_TC_OP_groupi_n_34 );
  assign csa_tree_ADD_TC_OP_groupi_n_42 = ~(csa_tree_ADD_TC_OP_groupi_n_29  ^ csa_tree_ADD_TC_OP_groupi_n_32 );
  assign csa_tree_ADD_TC_OP_groupi_n_41 = ~(csa_tree_ADD_TC_OP_groupi_n_20  | csa_tree_ADD_TC_OP_groupi_n_36 );
  assign csa_tree_ADD_TC_OP_groupi_n_40 = csa_tree_ADD_TC_OP_groupi_n_27  & csa_tree_ADD_TC_OP_groupi_n_37 ;
  assign csa_tree_ADD_TC_OP_groupi_n_39 = csa_tree_ADD_TC_OP_groupi_n_21  | csa_tree_ADD_TC_OP_groupi_n_35 ;
  assign out1[0] = ~(csa_tree_ADD_TC_OP_groupi_n_16  ^ in3[0] );
  assign csa_tree_ADD_TC_OP_groupi_n_37 = ~(csa_tree_ADD_TC_OP_groupi_n_23  ^ in3[2] );
  assign csa_tree_ADD_TC_OP_groupi_n_35 = ~csa_tree_ADD_TC_OP_groupi_n_36 ;
  assign csa_tree_ADD_TC_OP_groupi_n_36 = ~(csa_tree_ADD_TC_OP_groupi_n_25  ^ in3[1] );
  assign csa_tree_ADD_TC_OP_groupi_n_34 = ~(csa_tree_ADD_TC_OP_groupi_n_17  ^ csa_tree_ADD_TC_OP_groupi_n_24 );
  assign csa_tree_ADD_TC_OP_groupi_n_33 = ~(csa_tree_ADD_TC_OP_groupi_n_15  ^ csa_tree_ADD_TC_OP_groupi_n_19 );
  assign csa_tree_ADD_TC_OP_groupi_n_32 = ~(csa_tree_ADD_TC_OP_groupi_n_13  ^ in3[3] );
  assign csa_tree_ADD_TC_OP_groupi_n_31 = csa_tree_ADD_TC_OP_groupi_n_10  | csa_tree_ADD_TC_OP_groupi_n_16 ;
  assign csa_tree_ADD_TC_OP_groupi_n_30 = in3[1]  & csa_tree_ADD_TC_OP_groupi_n_26 ;
  assign csa_tree_ADD_TC_OP_groupi_n_29 = csa_tree_ADD_TC_OP_groupi_n_6  | csa_tree_ADD_TC_OP_groupi_n_23 ;
  assign csa_tree_ADD_TC_OP_groupi_n_28 = ~(csa_tree_ADD_TC_OP_groupi_n_15  | csa_tree_ADD_TC_OP_groupi_n_19 );
  assign csa_tree_ADD_TC_OP_groupi_n_27 = csa_tree_ADD_TC_OP_groupi_n_14  | csa_tree_ADD_TC_OP_groupi_n_18 ;
  assign csa_tree_ADD_TC_OP_groupi_n_26 = ~csa_tree_ADD_TC_OP_groupi_n_25 ;
  assign csa_tree_ADD_TC_OP_groupi_n_25 = csa_tree_ADD_TC_OP_groupi_n_9  | csa_tree_ADD_TC_OP_groupi_n_3 ;
  assign csa_tree_ADD_TC_OP_groupi_n_24 = csa_tree_ADD_TC_OP_groupi_n_8  | csa_tree_ADD_TC_OP_groupi_n_5 ;
  assign csa_tree_ADD_TC_OP_groupi_n_23 = csa_tree_ADD_TC_OP_groupi_n_8  | csa_tree_ADD_TC_OP_groupi_n_3 ;
  assign csa_tree_ADD_TC_OP_groupi_n_22 = csa_tree_ADD_TC_OP_groupi_n_9  | csa_tree_ADD_TC_OP_groupi_n_7 ;
  assign csa_tree_ADD_TC_OP_groupi_n_20 = ~csa_tree_ADD_TC_OP_groupi_n_21 ;
  assign csa_tree_ADD_TC_OP_groupi_n_21 = csa_tree_ADD_TC_OP_groupi_n_4  | csa_tree_ADD_TC_OP_groupi_n_5 ;
  assign csa_tree_ADD_TC_OP_groupi_n_19 = ~csa_tree_ADD_TC_OP_groupi_n_18 ;
  assign csa_tree_ADD_TC_OP_groupi_n_18 = in1[1]  & in2[1] ;
  assign csa_tree_ADD_TC_OP_groupi_n_17 = csa_tree_ADD_TC_OP_groupi_n_4  | csa_tree_ADD_TC_OP_groupi_n_12 ;
  assign csa_tree_ADD_TC_OP_groupi_n_16 = csa_tree_ADD_TC_OP_groupi_n_4  | csa_tree_ADD_TC_OP_groupi_n_2 ;
  assign csa_tree_ADD_TC_OP_groupi_n_15 = ~csa_tree_ADD_TC_OP_groupi_n_14 ;
  assign csa_tree_ADD_TC_OP_groupi_n_14 = in1[0]  & in2[2] ;
  assign csa_tree_ADD_TC_OP_groupi_n_13 = csa_tree_ADD_TC_OP_groupi_n_11  | csa_tree_ADD_TC_OP_groupi_n_2 ;
  assign csa_tree_ADD_TC_OP_groupi_n_12 = ~in2[3] ;
  assign csa_tree_ADD_TC_OP_groupi_n_11 = ~in1[3] ;
  assign csa_tree_ADD_TC_OP_groupi_n_10 = ~in3[0] ;
  assign csa_tree_ADD_TC_OP_groupi_n_9 = ~in1[1] ;
  assign csa_tree_ADD_TC_OP_groupi_n_8 = ~in1[2] ;
  assign csa_tree_ADD_TC_OP_groupi_n_7 = ~in2[2] ;
  assign csa_tree_ADD_TC_OP_groupi_n_6 = ~in3[2] ;
  assign csa_tree_ADD_TC_OP_groupi_n_5 = ~in2[1] ;
  assign csa_tree_ADD_TC_OP_groupi_n_4 = ~in1[0] ;
  assign csa_tree_ADD_TC_OP_groupi_n_3 = ~in2[0] ;
  assign csa_tree_ADD_TC_OP_groupi_n_2 = ~csa_tree_ADD_TC_OP_groupi_n_1 ;
  assign csa_tree_ADD_TC_OP_groupi_n_1 = ~csa_tree_ADD_TC_OP_groupi_n_3 ;
  assign csa_tree_ADD_TC_OP_groupi_n_0 = csa_tree_ADD_TC_OP_groupi_n_30  ^ csa_tree_ADD_TC_OP_groupi_n_44 ;
endmodule
