module top(in1, in2, in3, out1);
  input [3:0] in1, in2, in3;
  output [3:0] out1;
  wire [3:0] in1, in2, in3;
  wire [3:0] out1;
  wire csa_tree_ADD_TC_OP_1_groupi_n_0, csa_tree_ADD_TC_OP_1_groupi_n_1, csa_tree_ADD_TC_OP_1_groupi_n_2, csa_tree_ADD_TC_OP_1_groupi_n_3, csa_tree_ADD_TC_OP_1_groupi_n_4, csa_tree_ADD_TC_OP_1_groupi_n_5, csa_tree_ADD_TC_OP_1_groupi_n_6, csa_tree_ADD_TC_OP_1_groupi_n_7;
  wire csa_tree_ADD_TC_OP_1_groupi_n_8, csa_tree_ADD_TC_OP_1_groupi_n_9, csa_tree_ADD_TC_OP_1_groupi_n_10, csa_tree_ADD_TC_OP_1_groupi_n_11, csa_tree_ADD_TC_OP_1_groupi_n_12, csa_tree_ADD_TC_OP_1_groupi_n_13, csa_tree_ADD_TC_OP_1_groupi_n_14, csa_tree_ADD_TC_OP_1_groupi_n_15;
  wire csa_tree_ADD_TC_OP_1_groupi_n_16, csa_tree_ADD_TC_OP_1_groupi_n_17, csa_tree_ADD_TC_OP_1_groupi_n_18, csa_tree_ADD_TC_OP_1_groupi_n_19, csa_tree_ADD_TC_OP_1_groupi_n_21, csa_tree_ADD_TC_OP_1_groupi_n_22, csa_tree_ADD_TC_OP_1_groupi_n_23, csa_tree_ADD_TC_OP_1_groupi_n_24;
  wire csa_tree_ADD_TC_OP_1_groupi_n_25, csa_tree_ADD_TC_OP_1_groupi_n_26, csa_tree_ADD_TC_OP_1_groupi_n_27, csa_tree_ADD_TC_OP_1_groupi_n_29, csa_tree_ADD_TC_OP_1_groupi_n_30, csa_tree_ADD_TC_OP_1_groupi_n_31, csa_tree_ADD_TC_OP_1_groupi_n_32;
  assign out1[3] = ~(csa_tree_ADD_TC_OP_1_groupi_n_29  ^ csa_tree_ADD_TC_OP_1_groupi_n_32 );
  assign out1[2] = csa_tree_ADD_TC_OP_1_groupi_n_26  ^ csa_tree_ADD_TC_OP_1_groupi_n_30 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_32 = csa_tree_ADD_TC_OP_1_groupi_n_25  | csa_tree_ADD_TC_OP_1_groupi_n_31 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_31 = csa_tree_ADD_TC_OP_1_groupi_n_27  & csa_tree_ADD_TC_OP_1_groupi_n_26 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_30 = ~(csa_tree_ADD_TC_OP_1_groupi_n_5  ^ csa_tree_ADD_TC_OP_1_groupi_n_22 );
  assign csa_tree_ADD_TC_OP_1_groupi_n_29 = ~(csa_tree_ADD_TC_OP_1_groupi_n_17  ^ csa_tree_ADD_TC_OP_1_groupi_n_23 );
  assign out1[1] = csa_tree_ADD_TC_OP_1_groupi_n_16  ^ csa_tree_ADD_TC_OP_1_groupi_n_21 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_27 = csa_tree_ADD_TC_OP_1_groupi_n_6  | csa_tree_ADD_TC_OP_1_groupi_n_22 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_26 = csa_tree_ADD_TC_OP_1_groupi_n_19  | csa_tree_ADD_TC_OP_1_groupi_n_24 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_25 = csa_tree_ADD_TC_OP_1_groupi_n_6  & csa_tree_ADD_TC_OP_1_groupi_n_22 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_24 = csa_tree_ADD_TC_OP_1_groupi_n_16  & csa_tree_ADD_TC_OP_1_groupi_n_18 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_23 = ~(csa_tree_ADD_TC_OP_1_groupi_n_10  ^ in1[3] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_22 = ~(csa_tree_ADD_TC_OP_1_groupi_n_9  ^ in1[2] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_21 = ~(csa_tree_ADD_TC_OP_1_groupi_n_12  ^ in2[1] );
  assign out1[0] = ~(csa_tree_ADD_TC_OP_1_groupi_n_13  ^ in3[0] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_19 = ~(csa_tree_ADD_TC_OP_1_groupi_n_1  | csa_tree_ADD_TC_OP_1_groupi_n_12 );
  assign csa_tree_ADD_TC_OP_1_groupi_n_18 = in2[1]  | csa_tree_ADD_TC_OP_1_groupi_n_11 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_17 = csa_tree_ADD_TC_OP_1_groupi_n_7  | csa_tree_ADD_TC_OP_1_groupi_n_15 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_16 = csa_tree_ADD_TC_OP_1_groupi_n_4  | csa_tree_ADD_TC_OP_1_groupi_n_14 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_15 = in3[2]  & csa_tree_ADD_TC_OP_1_groupi_n_8 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_14 = in1[0]  & csa_tree_ADD_TC_OP_1_groupi_n_3 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_13 = ~(in1[0]  ^ in2[0] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_11 = ~csa_tree_ADD_TC_OP_1_groupi_n_12 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_12 = ~(in3[1]  ^ in1[1] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_10 = ~(in3[3]  ^ in2[3] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_9 = ~(in3[2]  ^ in2[2] );
  assign csa_tree_ADD_TC_OP_1_groupi_n_8 = in1[2]  | in2[2] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_7 = in1[2]  & in2[2] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_6 = ~csa_tree_ADD_TC_OP_1_groupi_n_5 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_5 = csa_tree_ADD_TC_OP_1_groupi_n_0  | csa_tree_ADD_TC_OP_1_groupi_n_2 ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_4 = in3[0]  & in2[0] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_3 = in3[0]  | in2[0] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_2 = ~in1[1] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_1 = ~in2[1] ;
  assign csa_tree_ADD_TC_OP_1_groupi_n_0 = ~in3[1] ;
endmodule
